module testbench();
// Declare inputs as regs and outputs as wires
reg clk;
reg [2:0] rs1;
reg [2:0] rs2;
reg [2:0] rd;
reg [7:0] write_data;
reg reg_write;
reg label_write;
reg label_read;

wire [7:0] regA_o;
wire [7:0] regB_o;

// Initialize all variables
initial begin        
	clk = 1;       // initial value of clock
	reg_write = 0;  	// initial value of reg_write
	label_write = 1;     // initial value of label_write
	label_read = 0;     // initial value of lable_read
	write_data = 8'b00000001;
	rs1 = 3'b001;
	rs2 = 3'b010;
	rd = 3'b001;

	#10  rd = 3'b010;
	write_data = 8'b10;
	#10  label_write = 0;
	reg_write = 1;
	write_data = 8'b11;
	#10  rd = 3'b001;
	write_data = 8'b100;
	#10  reg_write = 0;
	label_read = 1;
	write_data = 8'b101;
	

 end

// Clock generator
always begin
   #5  clk = ~clk; // Toggle clock every 5 ticks
						// this makes the clock cycle 10 ticks
end

// the following creates an instance of our program_counter register.
//   I copied this code verbatim from the walkthough.v that was
//   generated by Quartus when I created the .v file from the .bdf.

register_file	b2v_inst(
	.clk(clk),
	.reg_write(reg_write),
	.label_write(label_write),
	.label_read(label_read),
	.rd(rd),
	.rs1(rs1),
	.rs2(rs2),
	.write_data(write_data),
	.regA_o(regA_o),
	.regB_o(regB_o));



endmodule
